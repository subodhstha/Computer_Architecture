module and_gate (a, b, c);
    input a, b;
    output c;
    and and1(c, a, b);
endmodule