module or_gate (a, b, c);// module module_name(input, output)
    input a, b;
    output c;
    or or1(c, a, b);
endmodule